`timescale 1ns / 1ps

//
// This version of S-blocks does not generate warnings.
//
module SP_v2(
	input [47:0] din,
	output [31:0] dout
	);
	
// script generated
	wire [5:0] k0 = { din[0], din[5], din[1], din[2], din[3], din[4] };

	wire [3:0] S0 =
		k0 == 6'd0 ? 4'd14 :
		k0 == 6'd1 ? 4'd4 :
		k0 == 6'd2 ? 4'd13 :
		k0 == 6'd3 ? 4'd1 :
		k0 == 6'd4 ? 4'd2 :
		k0 == 6'd5 ? 4'd15 :
		k0 == 6'd6 ? 4'd11 :
		k0 == 6'd7 ? 4'd8 :
		k0 == 6'd8 ? 4'd3 :
		k0 == 6'd9 ? 4'd10 :
		k0 == 6'd10 ? 4'd6 :
		k0 == 6'd11 ? 4'd12 :
		k0 == 6'd12 ? 4'd5 :
		k0 == 6'd13 ? 4'd9 :
		k0 == 6'd14 ? 4'd0 :
		k0 == 6'd15 ? 4'd7 :

		k0 == 6'd16 ? 4'd0 :
		k0 == 6'd17 ? 4'd15 :
		k0 == 6'd18 ? 4'd7 :
		k0 == 6'd19 ? 4'd4 :
		k0 == 6'd20 ? 4'd14 :
		k0 == 6'd21 ? 4'd2 :
		k0 == 6'd22 ? 4'd13 :
		k0 == 6'd23 ? 4'd1 :
		k0 == 6'd24 ? 4'd10 :
		k0 == 6'd25 ? 4'd6 :
		k0 == 6'd26 ? 4'd12 :
		k0 == 6'd27 ? 4'd11 :
		k0 == 6'd28 ? 4'd9 :
		k0 == 6'd29 ? 4'd5 :
		k0 == 6'd30 ? 4'd3 :
		k0 == 6'd31 ? 4'd8 :

		k0 == 6'd32 ? 4'd4 :
		k0 == 6'd33 ? 4'd1 :
		k0 == 6'd34 ? 4'd14 :
		k0 == 6'd35 ? 4'd8 :
		k0 == 6'd36 ? 4'd13 :
		k0 == 6'd37 ? 4'd6 :
		k0 == 6'd38 ? 4'd2 :
		k0 == 6'd39 ? 4'd11 :
		k0 == 6'd40 ? 4'd15 :
		k0 == 6'd41 ? 4'd12 :
		k0 == 6'd42 ? 4'd9 :
		k0 == 6'd43 ? 4'd7 :
		k0 == 6'd44 ? 4'd3 :
		k0 == 6'd45 ? 4'd10 :
		k0 == 6'd46 ? 4'd5 :
		k0 == 6'd47 ? 4'd0 :

		k0 == 6'd48 ? 4'd15 :
		k0 == 6'd49 ? 4'd12 :
		k0 == 6'd50 ? 4'd8 :
		k0 == 6'd51 ? 4'd2 :
		k0 == 6'd52 ? 4'd4 :
		k0 == 6'd53 ? 4'd9 :
		k0 == 6'd54 ? 4'd1 :
		k0 == 6'd55 ? 4'd7 :
		k0 == 6'd56 ? 4'd5 :
		k0 == 6'd57 ? 4'd11 :
		k0 == 6'd58 ? 4'd3 :
		k0 == 6'd59 ? 4'd14 :
		k0 == 6'd60 ? 4'd10 :
		k0 == 6'd61 ? 4'd0 :
		k0 == 6'd62 ? 4'd6 :
		4'd13;

	wire [5:0] k1 = { din[6], din[11], din[7], din[8], din[9], din[10] };

	wire [3:0] S1 =
		k1 == 6'd0 ? 4'd15 :
		k1 == 6'd1 ? 4'd1 :
		k1 == 6'd2 ? 4'd8 :
		k1 == 6'd3 ? 4'd14 :
		k1 == 6'd4 ? 4'd6 :
		k1 == 6'd5 ? 4'd11 :
		k1 == 6'd6 ? 4'd3 :
		k1 == 6'd7 ? 4'd4 :
		k1 == 6'd8 ? 4'd9 :
		k1 == 6'd9 ? 4'd7 :
		k1 == 6'd10 ? 4'd2 :
		k1 == 6'd11 ? 4'd13 :
		k1 == 6'd12 ? 4'd12 :
		k1 == 6'd13 ? 4'd0 :
		k1 == 6'd14 ? 4'd5 :
		k1 == 6'd15 ? 4'd10 :

		k1 == 6'd16 ? 4'd3 :
		k1 == 6'd17 ? 4'd13 :
		k1 == 6'd18 ? 4'd4 :
		k1 == 6'd19 ? 4'd7 :
		k1 == 6'd20 ? 4'd15 :
		k1 == 6'd21 ? 4'd2 :
		k1 == 6'd22 ? 4'd8 :
		k1 == 6'd23 ? 4'd14 :
		k1 == 6'd24 ? 4'd12 :
		k1 == 6'd25 ? 4'd0 :
		k1 == 6'd26 ? 4'd1 :
		k1 == 6'd27 ? 4'd10 :
		k1 == 6'd28 ? 4'd6 :
		k1 == 6'd29 ? 4'd9 :
		k1 == 6'd30 ? 4'd11 :
		k1 == 6'd31 ? 4'd5 :

		k1 == 6'd32 ? 4'd0 :
		k1 == 6'd33 ? 4'd14 :
		k1 == 6'd34 ? 4'd7 :
		k1 == 6'd35 ? 4'd11 :
		k1 == 6'd36 ? 4'd10 :
		k1 == 6'd37 ? 4'd4 :
		k1 == 6'd38 ? 4'd13 :
		k1 == 6'd39 ? 4'd1 :
		k1 == 6'd40 ? 4'd5 :
		k1 == 6'd41 ? 4'd8 :
		k1 == 6'd42 ? 4'd12 :
		k1 == 6'd43 ? 4'd6 :
		k1 == 6'd44 ? 4'd9 :
		k1 == 6'd45 ? 4'd3 :
		k1 == 6'd46 ? 4'd2 :
		k1 == 6'd47 ? 4'd15 :

		k1 == 6'd48 ? 4'd13 :
		k1 == 6'd49 ? 4'd8 :
		k1 == 6'd50 ? 4'd10 :
		k1 == 6'd51 ? 4'd1 :
		k1 == 6'd52 ? 4'd3 :
		k1 == 6'd53 ? 4'd15 :
		k1 == 6'd54 ? 4'd4 :
		k1 == 6'd55 ? 4'd2 :
		k1 == 6'd56 ? 4'd11 :
		k1 == 6'd57 ? 4'd6 :
		k1 == 6'd58 ? 4'd7 :
		k1 == 6'd59 ? 4'd12 :
		k1 == 6'd60 ? 4'd0 :
		k1 == 6'd61 ? 4'd5 :
		k1 == 6'd62 ? 4'd14 :
		4'd9;

	wire [5:0] k2 = { din[12], din[17], din[13], din[14], din[15], din[16] };

	wire [3:0] S2 =
		k2 == 6'd0 ? 4'd10 :
		k2 == 6'd1 ? 4'd0 :
		k2 == 6'd2 ? 4'd9 :
		k2 == 6'd3 ? 4'd14 :
		k2 == 6'd4 ? 4'd6 :
		k2 == 6'd5 ? 4'd3 :
		k2 == 6'd6 ? 4'd15 :
		k2 == 6'd7 ? 4'd5 :
		k2 == 6'd8 ? 4'd1 :
		k2 == 6'd9 ? 4'd13 :
		k2 == 6'd10 ? 4'd12 :
		k2 == 6'd11 ? 4'd7 :
		k2 == 6'd12 ? 4'd11 :
		k2 == 6'd13 ? 4'd4 :
		k2 == 6'd14 ? 4'd2 :
		k2 == 6'd15 ? 4'd8 :

		k2 == 6'd16 ? 4'd13 :
		k2 == 6'd17 ? 4'd7 :
		k2 == 6'd18 ? 4'd0 :
		k2 == 6'd19 ? 4'd9 :
		k2 == 6'd20 ? 4'd3 :
		k2 == 6'd21 ? 4'd4 :
		k2 == 6'd22 ? 4'd6 :
		k2 == 6'd23 ? 4'd10 :
		k2 == 6'd24 ? 4'd2 :
		k2 == 6'd25 ? 4'd8 :
		k2 == 6'd26 ? 4'd5 :
		k2 == 6'd27 ? 4'd14 :
		k2 == 6'd28 ? 4'd12 :
		k2 == 6'd29 ? 4'd11 :
		k2 == 6'd30 ? 4'd15 :
		k2 == 6'd31 ? 4'd1 :

		k2 == 6'd32 ? 4'd13 :
		k2 == 6'd33 ? 4'd6 :
		k2 == 6'd34 ? 4'd4 :
		k2 == 6'd35 ? 4'd9 :
		k2 == 6'd36 ? 4'd8 :
		k2 == 6'd37 ? 4'd15 :
		k2 == 6'd38 ? 4'd3 :
		k2 == 6'd39 ? 4'd0 :
		k2 == 6'd40 ? 4'd11 :
		k2 == 6'd41 ? 4'd1 :
		k2 == 6'd42 ? 4'd2 :
		k2 == 6'd43 ? 4'd12 :
		k2 == 6'd44 ? 4'd5 :
		k2 == 6'd45 ? 4'd10 :
		k2 == 6'd46 ? 4'd14 :
		k2 == 6'd47 ? 4'd7 :

		k2 == 6'd48 ? 4'd1 :
		k2 == 6'd49 ? 4'd10 :
		k2 == 6'd50 ? 4'd13 :
		k2 == 6'd51 ? 4'd0 :
		k2 == 6'd52 ? 4'd6 :
		k2 == 6'd53 ? 4'd9 :
		k2 == 6'd54 ? 4'd8 :
		k2 == 6'd55 ? 4'd7 :
		k2 == 6'd56 ? 4'd4 :
		k2 == 6'd57 ? 4'd15 :
		k2 == 6'd58 ? 4'd14 :
		k2 == 6'd59 ? 4'd3 :
		k2 == 6'd60 ? 4'd11 :
		k2 == 6'd61 ? 4'd5 :
		k2 == 6'd62 ? 4'd2 :
		4'd12;

	wire [5:0] k3 = { din[18], din[23], din[19], din[20], din[21], din[22] };

	wire [3:0] S3 =
		k3 == 6'd0 ? 4'd7 :
		k3 == 6'd1 ? 4'd13 :
		k3 == 6'd2 ? 4'd14 :
		k3 == 6'd3 ? 4'd3 :
		k3 == 6'd4 ? 4'd0 :
		k3 == 6'd5 ? 4'd6 :
		k3 == 6'd6 ? 4'd9 :
		k3 == 6'd7 ? 4'd10 :
		k3 == 6'd8 ? 4'd1 :
		k3 == 6'd9 ? 4'd2 :
		k3 == 6'd10 ? 4'd8 :
		k3 == 6'd11 ? 4'd5 :
		k3 == 6'd12 ? 4'd11 :
		k3 == 6'd13 ? 4'd12 :
		k3 == 6'd14 ? 4'd4 :
		k3 == 6'd15 ? 4'd15 :

		k3 == 6'd16 ? 4'd13 :
		k3 == 6'd17 ? 4'd8 :
		k3 == 6'd18 ? 4'd11 :
		k3 == 6'd19 ? 4'd5 :
		k3 == 6'd20 ? 4'd6 :
		k3 == 6'd21 ? 4'd15 :
		k3 == 6'd22 ? 4'd0 :
		k3 == 6'd23 ? 4'd3 :
		k3 == 6'd24 ? 4'd4 :
		k3 == 6'd25 ? 4'd7 :
		k3 == 6'd26 ? 4'd2 :
		k3 == 6'd27 ? 4'd12 :
		k3 == 6'd28 ? 4'd1 :
		k3 == 6'd29 ? 4'd10 :
		k3 == 6'd30 ? 4'd14 :
		k3 == 6'd31 ? 4'd9 :

		k3 == 6'd32 ? 4'd10 :
		k3 == 6'd33 ? 4'd6 :
		k3 == 6'd34 ? 4'd9 :
		k3 == 6'd35 ? 4'd0 :
		k3 == 6'd36 ? 4'd12 :
		k3 == 6'd37 ? 4'd11 :
		k3 == 6'd38 ? 4'd7 :
		k3 == 6'd39 ? 4'd13 :
		k3 == 6'd40 ? 4'd15 :
		k3 == 6'd41 ? 4'd1 :
		k3 == 6'd42 ? 4'd3 :
		k3 == 6'd43 ? 4'd14 :
		k3 == 6'd44 ? 4'd5 :
		k3 == 6'd45 ? 4'd2 :
		k3 == 6'd46 ? 4'd8 :
		k3 == 6'd47 ? 4'd4 :

		k3 == 6'd48 ? 4'd3 :
		k3 == 6'd49 ? 4'd15 :
		k3 == 6'd50 ? 4'd0 :
		k3 == 6'd51 ? 4'd6 :
		k3 == 6'd52 ? 4'd10 :
		k3 == 6'd53 ? 4'd1 :
		k3 == 6'd54 ? 4'd13 :
		k3 == 6'd55 ? 4'd8 :
		k3 == 6'd56 ? 4'd9 :
		k3 == 6'd57 ? 4'd4 :
		k3 == 6'd58 ? 4'd5 :
		k3 == 6'd59 ? 4'd11 :
		k3 == 6'd60 ? 4'd12 :
		k3 == 6'd61 ? 4'd7 :
		k3 == 6'd62 ? 4'd2 :
		4'd14;

	wire [5:0] k4 = { din[24], din[29], din[25], din[26], din[27], din[28] };

	wire [3:0] S4 =
		k4 == 6'd0 ? 4'd2 :
		k4 == 6'd1 ? 4'd12 :
		k4 == 6'd2 ? 4'd4 :
		k4 == 6'd3 ? 4'd1 :
		k4 == 6'd4 ? 4'd7 :
		k4 == 6'd5 ? 4'd10 :
		k4 == 6'd6 ? 4'd11 :
		k4 == 6'd7 ? 4'd6 :
		k4 == 6'd8 ? 4'd8 :
		k4 == 6'd9 ? 4'd5 :
		k4 == 6'd10 ? 4'd3 :
		k4 == 6'd11 ? 4'd15 :
		k4 == 6'd12 ? 4'd13 :
		k4 == 6'd13 ? 4'd0 :
		k4 == 6'd14 ? 4'd14 :
		k4 == 6'd15 ? 4'd9 :

		k4 == 6'd16 ? 4'd14 :
		k4 == 6'd17 ? 4'd11 :
		k4 == 6'd18 ? 4'd2 :
		k4 == 6'd19 ? 4'd12 :
		k4 == 6'd20 ? 4'd4 :
		k4 == 6'd21 ? 4'd7 :
		k4 == 6'd22 ? 4'd13 :
		k4 == 6'd23 ? 4'd1 :
		k4 == 6'd24 ? 4'd5 :
		k4 == 6'd25 ? 4'd0 :
		k4 == 6'd26 ? 4'd15 :
		k4 == 6'd27 ? 4'd10 :
		k4 == 6'd28 ? 4'd3 :
		k4 == 6'd29 ? 4'd9 :
		k4 == 6'd30 ? 4'd8 :
		k4 == 6'd31 ? 4'd6 :

		k4 == 6'd32 ? 4'd4 :
		k4 == 6'd33 ? 4'd2 :
		k4 == 6'd34 ? 4'd1 :
		k4 == 6'd35 ? 4'd11 :
		k4 == 6'd36 ? 4'd10 :
		k4 == 6'd37 ? 4'd13 :
		k4 == 6'd38 ? 4'd7 :
		k4 == 6'd39 ? 4'd8 :
		k4 == 6'd40 ? 4'd15 :
		k4 == 6'd41 ? 4'd9 :
		k4 == 6'd42 ? 4'd12 :
		k4 == 6'd43 ? 4'd5 :
		k4 == 6'd44 ? 4'd6 :
		k4 == 6'd45 ? 4'd3 :
		k4 == 6'd46 ? 4'd0 :
		k4 == 6'd47 ? 4'd14 :

		k4 == 6'd48 ? 4'd11 :
		k4 == 6'd49 ? 4'd8 :
		k4 == 6'd50 ? 4'd12 :
		k4 == 6'd51 ? 4'd7 :
		k4 == 6'd52 ? 4'd1 :
		k4 == 6'd53 ? 4'd14 :
		k4 == 6'd54 ? 4'd2 :
		k4 == 6'd55 ? 4'd13 :
		k4 == 6'd56 ? 4'd6 :
		k4 == 6'd57 ? 4'd15 :
		k4 == 6'd58 ? 4'd0 :
		k4 == 6'd59 ? 4'd9 :
		k4 == 6'd60 ? 4'd10 :
		k4 == 6'd61 ? 4'd4 :
		k4 == 6'd62 ? 4'd5 :
		4'd3;

	wire [5:0] k5 = { din[30], din[35], din[31], din[32], din[33], din[34] };

	wire [3:0] S5 =
		k5 == 6'd0 ? 4'd12 :
		k5 == 6'd1 ? 4'd1 :
		k5 == 6'd2 ? 4'd10 :
		k5 == 6'd3 ? 4'd15 :
		k5 == 6'd4 ? 4'd9 :
		k5 == 6'd5 ? 4'd2 :
		k5 == 6'd6 ? 4'd6 :
		k5 == 6'd7 ? 4'd8 :
		k5 == 6'd8 ? 4'd0 :
		k5 == 6'd9 ? 4'd13 :
		k5 == 6'd10 ? 4'd3 :
		k5 == 6'd11 ? 4'd4 :
		k5 == 6'd12 ? 4'd14 :
		k5 == 6'd13 ? 4'd7 :
		k5 == 6'd14 ? 4'd5 :
		k5 == 6'd15 ? 4'd11 :

		k5 == 6'd16 ? 4'd10 :
		k5 == 6'd17 ? 4'd15 :
		k5 == 6'd18 ? 4'd4 :
		k5 == 6'd19 ? 4'd2 :
		k5 == 6'd20 ? 4'd7 :
		k5 == 6'd21 ? 4'd12 :
		k5 == 6'd22 ? 4'd9 :
		k5 == 6'd23 ? 4'd5 :
		k5 == 6'd24 ? 4'd6 :
		k5 == 6'd25 ? 4'd1 :
		k5 == 6'd26 ? 4'd13 :
		k5 == 6'd27 ? 4'd14 :
		k5 == 6'd28 ? 4'd0 :
		k5 == 6'd29 ? 4'd11 :
		k5 == 6'd30 ? 4'd3 :
		k5 == 6'd31 ? 4'd8 :

		k5 == 6'd32 ? 4'd9 :
		k5 == 6'd33 ? 4'd14 :
		k5 == 6'd34 ? 4'd15 :
		k5 == 6'd35 ? 4'd5 :
		k5 == 6'd36 ? 4'd2 :
		k5 == 6'd37 ? 4'd8 :
		k5 == 6'd38 ? 4'd12 :
		k5 == 6'd39 ? 4'd3 :
		k5 == 6'd40 ? 4'd7 :
		k5 == 6'd41 ? 4'd0 :
		k5 == 6'd42 ? 4'd4 :
		k5 == 6'd43 ? 4'd10 :
		k5 == 6'd44 ? 4'd1 :
		k5 == 6'd45 ? 4'd13 :
		k5 == 6'd46 ? 4'd11 :
		k5 == 6'd47 ? 4'd6 :

		k5 == 6'd48 ? 4'd4 :
		k5 == 6'd49 ? 4'd3 :
		k5 == 6'd50 ? 4'd2 :
		k5 == 6'd51 ? 4'd12 :
		k5 == 6'd52 ? 4'd9 :
		k5 == 6'd53 ? 4'd5 :
		k5 == 6'd54 ? 4'd15 :
		k5 == 6'd55 ? 4'd10 :
		k5 == 6'd56 ? 4'd11 :
		k5 == 6'd57 ? 4'd14 :
		k5 == 6'd58 ? 4'd1 :
		k5 == 6'd59 ? 4'd7 :
		k5 == 6'd60 ? 4'd6 :
		k5 == 6'd61 ? 4'd0 :
		k5 == 6'd62 ? 4'd8 :
		4'd13;

	wire [5:0] k6 = { din[36], din[41], din[37], din[38], din[39], din[40] };

	wire [3:0] S6 =
		k6 == 6'd0 ? 4'd4 :
		k6 == 6'd1 ? 4'd11 :
		k6 == 6'd2 ? 4'd2 :
		k6 == 6'd3 ? 4'd14 :
		k6 == 6'd4 ? 4'd15 :
		k6 == 6'd5 ? 4'd0 :
		k6 == 6'd6 ? 4'd8 :
		k6 == 6'd7 ? 4'd13 :
		k6 == 6'd8 ? 4'd3 :
		k6 == 6'd9 ? 4'd12 :
		k6 == 6'd10 ? 4'd9 :
		k6 == 6'd11 ? 4'd7 :
		k6 == 6'd12 ? 4'd5 :
		k6 == 6'd13 ? 4'd10 :
		k6 == 6'd14 ? 4'd6 :
		k6 == 6'd15 ? 4'd1 :

		k6 == 6'd16 ? 4'd13 :
		k6 == 6'd17 ? 4'd0 :
		k6 == 6'd18 ? 4'd11 :
		k6 == 6'd19 ? 4'd7 :
		k6 == 6'd20 ? 4'd4 :
		k6 == 6'd21 ? 4'd9 :
		k6 == 6'd22 ? 4'd1 :
		k6 == 6'd23 ? 4'd10 :
		k6 == 6'd24 ? 4'd14 :
		k6 == 6'd25 ? 4'd3 :
		k6 == 6'd26 ? 4'd5 :
		k6 == 6'd27 ? 4'd12 :
		k6 == 6'd28 ? 4'd2 :
		k6 == 6'd29 ? 4'd15 :
		k6 == 6'd30 ? 4'd8 :
		k6 == 6'd31 ? 4'd6 :

		k6 == 6'd32 ? 4'd1 :
		k6 == 6'd33 ? 4'd4 :
		k6 == 6'd34 ? 4'd11 :
		k6 == 6'd35 ? 4'd13 :
		k6 == 6'd36 ? 4'd12 :
		k6 == 6'd37 ? 4'd3 :
		k6 == 6'd38 ? 4'd7 :
		k6 == 6'd39 ? 4'd14 :
		k6 == 6'd40 ? 4'd10 :
		k6 == 6'd41 ? 4'd15 :
		k6 == 6'd42 ? 4'd6 :
		k6 == 6'd43 ? 4'd8 :
		k6 == 6'd44 ? 4'd0 :
		k6 == 6'd45 ? 4'd5 :
		k6 == 6'd46 ? 4'd9 :
		k6 == 6'd47 ? 4'd2 :

		k6 == 6'd48 ? 4'd6 :
		k6 == 6'd49 ? 4'd11 :
		k6 == 6'd50 ? 4'd13 :
		k6 == 6'd51 ? 4'd8 :
		k6 == 6'd52 ? 4'd1 :
		k6 == 6'd53 ? 4'd4 :
		k6 == 6'd54 ? 4'd10 :
		k6 == 6'd55 ? 4'd7 :
		k6 == 6'd56 ? 4'd9 :
		k6 == 6'd57 ? 4'd5 :
		k6 == 6'd58 ? 4'd0 :
		k6 == 6'd59 ? 4'd15 :
		k6 == 6'd60 ? 4'd14 :
		k6 == 6'd61 ? 4'd2 :
		k6 == 6'd62 ? 4'd3 :
		4'd12;

	wire [5:0] k7 = { din[42], din[47], din[43], din[44], din[45], din[46] };

	wire [3:0] S7 =
		k7 == 6'd0 ? 4'd13 :
		k7 == 6'd1 ? 4'd2 :
		k7 == 6'd2 ? 4'd8 :
		k7 == 6'd3 ? 4'd4 :
		k7 == 6'd4 ? 4'd6 :
		k7 == 6'd5 ? 4'd15 :
		k7 == 6'd6 ? 4'd11 :
		k7 == 6'd7 ? 4'd1 :
		k7 == 6'd8 ? 4'd10 :
		k7 == 6'd9 ? 4'd9 :
		k7 == 6'd10 ? 4'd3 :
		k7 == 6'd11 ? 4'd14 :
		k7 == 6'd12 ? 4'd5 :
		k7 == 6'd13 ? 4'd0 :
		k7 == 6'd14 ? 4'd12 :
		k7 == 6'd15 ? 4'd7 :

		k7 == 6'd16 ? 4'd1 :
		k7 == 6'd17 ? 4'd15 :
		k7 == 6'd18 ? 4'd13 :
		k7 == 6'd19 ? 4'd8 :
		k7 == 6'd20 ? 4'd10 :
		k7 == 6'd21 ? 4'd3 :
		k7 == 6'd22 ? 4'd7 :
		k7 == 6'd23 ? 4'd4 :
		k7 == 6'd24 ? 4'd12 :
		k7 == 6'd25 ? 4'd5 :
		k7 == 6'd26 ? 4'd6 :
		k7 == 6'd27 ? 4'd11 :
		k7 == 6'd28 ? 4'd0 :
		k7 == 6'd29 ? 4'd14 :
		k7 == 6'd30 ? 4'd9 :
		k7 == 6'd31 ? 4'd2 :

		k7 == 6'd32 ? 4'd7 :
		k7 == 6'd33 ? 4'd11 :
		k7 == 6'd34 ? 4'd4 :
		k7 == 6'd35 ? 4'd1 :
		k7 == 6'd36 ? 4'd9 :
		k7 == 6'd37 ? 4'd12 :
		k7 == 6'd38 ? 4'd14 :
		k7 == 6'd39 ? 4'd2 :
		k7 == 6'd40 ? 4'd0 :
		k7 == 6'd41 ? 4'd6 :
		k7 == 6'd42 ? 4'd10 :
		k7 == 6'd43 ? 4'd13 :
		k7 == 6'd44 ? 4'd15 :
		k7 == 6'd45 ? 4'd3 :
		k7 == 6'd46 ? 4'd5 :
		k7 == 6'd47 ? 4'd8 :

		k7 == 6'd48 ? 4'd2 :
		k7 == 6'd49 ? 4'd1 :
		k7 == 6'd50 ? 4'd14 :
		k7 == 6'd51 ? 4'd7 :
		k7 == 6'd52 ? 4'd4 :
		k7 == 6'd53 ? 4'd10 :
		k7 == 6'd54 ? 4'd8 :
		k7 == 6'd55 ? 4'd13 :
		k7 == 6'd56 ? 4'd15 :
		k7 == 6'd57 ? 4'd12 :
		k7 == 6'd58 ? 4'd9 :
		k7 == 6'd59 ? 4'd0 :
		k7 == 6'd60 ? 4'd3 :
		k7 == 6'd61 ? 4'd5 :
		k7 == 6'd62 ? 4'd6 :
		4'd11;
// end script generated

	wire [31:0] dtmp = {
		S7[0], S7[1], S7[2], S7[3],
		S6[0], S6[1], S6[2], S6[3],
		S5[0], S5[1], S5[2], S5[3],
		S4[0], S4[1], S4[2], S4[3],
		S3[0], S3[1], S3[2], S3[3],
		S2[0], S2[1], S2[2], S2[3],
		S1[0], S1[1], S1[2], S1[3],
		S0[0], S0[1], S0[2], S0[3]
	};

	assign dout = {
		dtmp[24], dtmp[3], dtmp[10], dtmp[21], dtmp[5], dtmp[29], dtmp[12], dtmp[18], 
		dtmp[8], dtmp[2], dtmp[26], dtmp[31], dtmp[13], dtmp[23], dtmp[7], dtmp[1], 
		dtmp[9], dtmp[30], dtmp[17], dtmp[4], dtmp[25], dtmp[22], dtmp[14], dtmp[0], 
		dtmp[16], dtmp[27], dtmp[11], dtmp[28], dtmp[20], dtmp[19], dtmp[6], dtmp[15]
	};


endmodule
